module Smg(
    input wire [1:0]d_m,           // 显示距离费用，起步价和单价的选择信号，0表示显示单价起步价，1表示显示距离费用
    input wire [31:0] data_fx,    // 费用信号，16位
    input wire [31:0] data_tm,  // 距离信号，16位
	 input wire [31:0] data_zk,  // 起步价
    input wire [2:0] Bit_Sel,    // 数码管位选信号，3位
    output reg [7:0] Seg,    // 数码管段选信号，8位
    output reg [2:0] AN      // 数码管位选信号，2位
);
    reg [3:0] Data_now;      // 当前需要显示的数据
    initial 
    begin 
        Data_now = 4'b0;    // 初始化当前需要显示的数据为0
        Seg = 8'b0;   // 初始化数码管段选控制信号为0
    end
      
    always @(*)   // 根据位选信号控制数码管位选信号
    begin
        case(Bit_Sel)
            3'b000: AN<=3'b000;    // 选择第一位数码管
            3'b001: AN<=3'b001;    // 选择第二位数码管
            3'b010: AN<=3'b010;    // 选择第三位数码管
            3'b011: AN<=3'b011;    // 选择第四位数码管
				3'b100: AN<=3'b100;    // 选择第五位数码管
            3'b101: AN<=3'b101;    // 选择第六位数码管
            3'b110: AN<=3'b110;    // 选择第七位数码管
            3'b111: AN<=3'b111;    // 选择第八位数码管
            default: AN<=3'b111;  // 默认为不显示任何数码管
        endcase
    end
    
    always @(*)    // 根据显示距离还是费用的选择信号和位选信号，确定需要显示的数据
    begin
        if(d_m==2'b00)   // 如果选择显示距离费用，则从距离费用信号中选择需要显示的数据
        begin
            case(Bit_Sel)
                3'b000: Data_now[3:0] <= data_fx[31:28];   // 选择距离信号的高4位
                3'b001: Data_now[3:0] <= data_fx[27:24];    // 选择距离信号的第2~5位
                3'b010: Data_now[3:0] <= data_fx[23:20];     // 选择距离信号的第6~9位
                3'b011: Data_now[3:0] <= data_fx[19:16];     // 选择距离信号的低4位
					 3'b100: Data_now[3:0] <= data_fx[15:12];   // 选择距离信号的高4位
                3'b101: Data_now[3:0] <= data_fx[11:8];    // 选择距离信号的第2~5位
                3'b110: Data_now[3:0] <= data_fx[7:4];     // 选择距离信号的第6~9位
                3'b111: Data_now[3:0] <= data_fx[3:0];     // 选择距离信号的低4位
                default: Data_now[3:0] <= data_fx[31:28];   // 默认选择距离信号的低4位
            endcase
        end
        else if(d_m==2'b01)   // 如果选择显示启程价和单价，则从启程价和单价信号中选择需要显示的数据
        begin
			   case(Bit_Sel)
                3'b000: Data_now[3:0] <= data_tm[31:28];   // 选择距离信号的高4位
                3'b001: Data_now[3:0] <= data_tm[27:24];    // 选择距离信号的第2~5位
                3'b010: Data_now[3:0] <= data_tm[23:20];     // 选择距离信号的第6~9位
                3'b011: Data_now[3:0] <= data_tm[19:16];     // 选择距离信号的低4位
					 3'b100: Data_now[3:0] <= data_tm[15:12];   // 选择距离信号的高4位
                3'b101: Data_now[3:0] <= data_tm[11:8];    // 选择距离信号的第2~5位
                3'b110: Data_now[3:0] <= data_tm[7:4];     // 选择距离信号的第6~9位
                3'b111: Data_now[3:0] <= data_tm[3:0];     // 选择距离信号的低4位
                default: Data_now[3:0] <= data_tm[31:28];   // 默认选择距离信号的低4位
            endcase
		  end
		  else if(d_m==2'b10)   // 如果选择显示启程价和单价，则从启程价和单价信号中选择需要显示的数据
        begin
			   case(Bit_Sel)
                3'b000: Data_now[3:0] <= data_zk[31:28];   // 选择距离信号的高4位
                3'b001: Data_now[3:0] <= data_zk[27:24];    // 选择距离信号的第2~5位
                3'b010: Data_now[3:0] <= data_zk[23:20];     // 选择距离信号的第6~9位
                3'b011: Data_now[3:0] <= data_zk[19:16];     // 选择距离信号的低4位
					 3'b100: Data_now[3:0] <= data_zk[15:12];   // 选择距离信号的高4位
                3'b101: Data_now[3:0] <= data_zk[11:8];    // 选择距离信号的第2~5位
                3'b110: Data_now[3:0] <= data_zk[7:4];     // 选择距离信号的第6~9位
                3'b111: Data_now[3:0] <= data_zk[3:0];     // 选择距离信号的低4位
                default: Data_now[3:0] <= data_zk[31:28];   // 默认选择距离信号的低4位
            endcase
		  end
		   else  // 如果选择显示启程价和单价，则从启程价和单价信号中选择需要显示的数据
        begin
			   case(Bit_Sel)
                3'b000: Data_now[3:0] <= data_tm[31:28];   // 选择距离信号的高4位
                3'b001: Data_now[3:0] <= data_tm[27:24];    // 选择距离信号的第2~5位
                3'b010: Data_now[3:0] <= data_tm[23:20];     // 选择距离信号的第6~9位
                3'b011: Data_now[3:0] <= data_tm[19:16];     // 选择距离信号的低4位
					 3'b100: Data_now[3:0] <= data_tm[15:12];   // 选择距离信号的高4位
                3'b101: Data_now[3:0] <= data_tm[11:8];    // 选择距离信号的第2~5位
                3'b110: Data_now[3:0] <= data_tm[7:4];     // 选择距离信号的第6~9位
                3'b111: Data_now[3:0] <= data_tm[3:0];     // 选择距离信号的低4位
                default: Data_now[3:0] <= data_tm[31:28];   // 默认选择距离信号的低4位
            endcase
		  end
	 end
	 
	 always @(*)
	 begin
	  begin 
			// 根据 Data_now 的低 4 位数字选择对应的信号，点亮数码管
			case(Data_now[3:0])
				 // 数字 0 的信号
				 4'b0000: Seg[7:0] <= 8'b0011_1111;
				 // 数字 1 的信号
				 4'b0001: Seg[7:0] <= 8'b0000_0110;
				 // 数字 2 的信号
				 4'b0010: Seg[7:0] <= 8'b0101_1011;
				 // 数字 3 的信号
				 4'b0011: Seg[7:0] <= 8'b0100_1111;
				 // 数字 4 的信号
				 4'b0100: Seg[7:0] <= 8'b0110_0110;
				 // 数字 5 的信号
				 4'b0101: Seg[7:0] <= 8'b0110_1101;
				 // 数字 6 的信号
				 4'b0110: Seg[7:0] <= 8'b0111_1101;
				 // 数字 7 的信号
				 4'b0111: Seg[7:0] <= 8'b0000_0111;
				 // 数字 8 的信号
				 4'b1000: Seg[7:0] <= 8'b0111_1111;
				 // 数字 9 的信号
				 4'b1001: Seg[7:0] <= 8'b0110_1111;
				 // 其他数字不显示
				 default: Seg[7:0] <= 8'b0100_0000;  // .
			endcase
	  end   
    end

endmodule
